library verilog;
use verilog.vl_types.all;
entity counter10x4_vlg_tst is
end counter10x4_vlg_tst;
